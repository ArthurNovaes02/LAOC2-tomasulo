module FPmultipliers (Clock, CDB, )
  input Clock;
  output CDB;
end module
